// Copyright (C) 2024  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 23.1std.1 Build 993 05/14/2024 SC Standard Edition"
// CREATED		"Fri Feb 14 12:18:15 2025"

module counter(
	CLK,
	RST,
	count0,
	count1,
	count2,
	count3,
	count4,
	count5,
	count6,
	count7
);


input wire	CLK;
input wire	RST;
output wire	count0;
output wire	count1;
output wire	count2;
output wire	count3;
output wire	count4;
output wire	count5;
output wire	count6;
output wire	count7;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;

assign	count3 = SYNTHESIZED_WIRE_5;
assign	SYNTHESIZED_WIRE_2 = 1;
assign	SYNTHESIZED_WIRE_4 = 0;




four_bit_counter	b2v_inst(
	.clk(SYNTHESIZED_WIRE_0),
	.reset(RST),
	.count_0(count0),
	.count_1(count1),
	.count_2(count2),
	.count_3(SYNTHESIZED_WIRE_5));




four_bit_counter	b2v_inst3(
	.clk(SYNTHESIZED_WIRE_1),
	.reset(RST),
	.count_0(count4),
	.count_1(count5),
	.count_2(count6),
	.count_3(count7));

assign	SYNTHESIZED_WIRE_3 =  ~CLK;

assign	SYNTHESIZED_WIRE_0 = ~(SYNTHESIZED_WIRE_2 & SYNTHESIZED_WIRE_3);

assign	SYNTHESIZED_WIRE_6 =  ~SYNTHESIZED_WIRE_4;

assign	SYNTHESIZED_WIRE_1 = ~(SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_6);


endmodule
