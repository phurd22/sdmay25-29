// Copyright (C) 2024  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 23.1std.1 Build 993 05/14/2024 SC Standard Edition"
// CREATED		"Mon Mar 10 14:37:01 2025"

module addr_plus_one_4bit(
	decade_addr,
	rst_n,
	decade_1_addr
);


input wire	[3:0] decade_addr;
output wire	rst_n;
output wire	[3:0] decade_1_addr;

wire	[3:0] decade_1_addr_ALTERA_SYNTHESIZED;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_4;

assign	SYNTHESIZED_WIRE_6 = 0;
assign	SYNTHESIZED_WIRE_4 = 1;



assign	rst_n =  ~SYNTHESIZED_WIRE_0;




adder_4bit	b2v_inst5(
	.X3(decade_addr[3]),
	.Y3(SYNTHESIZED_WIRE_6),
	.X2(decade_addr[2]),
	.Y2(SYNTHESIZED_WIRE_6),
	.X1(decade_addr[1]),
	.Y1(SYNTHESIZED_WIRE_6),
	.X0(decade_addr[0]),
	.Y0(SYNTHESIZED_WIRE_4),
	.Ci(SYNTHESIZED_WIRE_6),
	.S0(decade_1_addr_ALTERA_SYNTHESIZED[0]),
	.S1(decade_1_addr_ALTERA_SYNTHESIZED[1]),
	.S2(decade_1_addr_ALTERA_SYNTHESIZED[2]),
	.S3(decade_1_addr_ALTERA_SYNTHESIZED[3]),
	.Co(SYNTHESIZED_WIRE_0));

assign	decade_1_addr = decade_1_addr_ALTERA_SYNTHESIZED;

endmodule
