// Copyright (C) 2024  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 23.1std.1 Build 993 05/14/2024 SC Standard Edition"
// CREATED		"Fri Feb 21 13:23:57 2025"

module HolderShifterModule(
	DCLK,
	shift1,
	RST,
	HS_Input,
	HS_Output
);

input wire	DCLK;
input wire	shift1;
input wire	RST;
input wire	HS_Input;
output wire	HS_Output;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
reg	DFF_inst;

assign	SYNTHESIZED_WIRE_1 = 1;

always@(posedge DCLK or negedge SYNTHESIZED_WIRE_0 or negedge SYNTHESIZED_WIRE_1)
begin
if (!SYNTHESIZED_WIRE_0)
	begin
	DFF_inst <= 0;
	end
else
if (!SYNTHESIZED_WIRE_1)
	begin
	DFF_inst <= 1;
	end
else
	begin
	DFF_inst <= HS_Input;
	end
end

assign	SYNTHESIZED_WIRE_0 =  ~RST;

// Instantiate the 2-to-1 multiplexer
TwotoOneMux b2v_inst5(
	.Zero(DFF_inst),
	.S(shift1),
	.One(HS_Input),
	.f(HS_Output));

endmodule

// 2-to-1 Multiplexer module definition
module TwotoOneMux(
    input wire Zero,     // Input 0
    input wire One,      // Input 1
    input wire S,        // Selector signal
    output wire f        // Output
);
    assign f = (S) ? One : Zero;
endmodule

