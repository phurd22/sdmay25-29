module sevens_eeprom (
    input wire clk,            // Clock signal
    input wire rst_n,          // Active-low reset
    input wire cs_n,           // Active-low chip select
    input wire oe_n,           // Active-low output enable
    input wire [15:0] addr,   // 16-bit address bus
    output wire [7:0] data    // 8-bit data bus (output only)
);

    // Memory size is fixed at 2^16 = 65,536 locations
    reg [7:0] memory [0:65535];

    // Initialize memory with hard-coded dummy data
	 initial begin
    memory[0] = 2'h01;
	 memory[1] = 2'h03;
	 memory[2] = 2'h07;
	 memory[3] = 2'h0c;
	 memory[4] = 2'h1c;
	 
	 memory[5] = 2'h34;
	 memory[6] = 2'h7a;
	 memory[7] = 2'hc4;
	 memory[8] = 2'hd8;
	 memory[9] = 2'h6c;
	 
	 memory[10] = 2'he0;
	 memory[11] = 2'he8;
	 memory[12] = 2'h98;
	 memory[13] = 2'h20;
	 memory[14] = 2'h40;
	 
	 memory[15] = 2'h60;
	 memory[16] = 2'h10;
	 memory[17] = 2'h60;
	 memory[18] = 2'h80;
	 memory[19] = 2'he0;
	 
	 memory[20] = 2'h00;
	 memory[21] = 2'hc0;
	 memory[22] = 2'h40;
	 memory[23] = 2'h00;
	 memory[24] = 2'h00;
	 
	 memory[25] = 2'h00;
	 memory[26] = 2'h00;
	 memory[27] = 2'h00;
	 memory[28] = 2'h00;
	 memory[29] = 2'h00;
	 
	 end

    // Internal data register
    reg [7:0] data_out;

    // Tri-state buffer control
    assign data = (!cs_n && !oe_n) ? data_out : 8'bz;

    // Read operation
    always @(*) begin
        if (!cs_n && !oe_n) begin
            // Read data from memory when output enable is active
            data_out = memory[addr];
        end else begin
            data_out = 8'bz;
        end
    end

endmodule